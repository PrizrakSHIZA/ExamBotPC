    ����          @ExamBotPC, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null   xSystem.Collections.Generic.List`1[[ExamTrainBot.User, ExamBotPC, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  ExamTrainBot.User[]   	                   ExamTrainBot.User   	      ExamTrainBot.User   idname
subscriberisadminontestcurrentquestiontestcreationpointscompletedtestsmistakesdate       	~System.Collections.Generic.List`1[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]~System.Collections.Generic.List`1[[ExamTrainBot.Tests.Test, ExamBotPC, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null]]�System.Collections.Generic.List`1[[System.Boolean[], mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   ��8=       Ефим Ряскин       	   	   	    @Ɖ��   ~System.Collections.Generic.List`1[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   _items_size_version  		            ~System.Collections.Generic.List`1[[ExamTrainBot.Tests.Test, ExamBotPC, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  ExamTrainBot.Tests.Test[]   	
            �System.Collections.Generic.List`1[[System.Boolean[], mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   _items_size_version  System.Boolean[][]	         	         
          ExamTrainBot.Tests.Test   	            	   


   ExamTrainBot.Tests.Test   Text	questions�System.Collections.Generic.List`1[[ExamTrainBot.Tests.Questions.Question, ExamBotPC, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null]]      New rule	               �System.Collections.Generic.List`1[[ExamTrainBot.Tests.Questions.Question, ExamBotPC, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  'ExamTrainBot.Tests.Questions.Question[]   	                   %ExamTrainBot.Tests.Questions.Question   	   	   	   
   )ExamTrainBot.Tests.Questions.TestQuestion   <text>k__BackingField<points>k__BackingField<variants>k__BackingFieldcolumns<answer>k__BackingField        Answer is 5   	         5   /ExamTrainBot.Tests.Questions.ConformityQuestion   <text>k__BackingField<points>k__BackingField<answer>k__BackingField<variants>k__BackingFieldruledelimiterChars       Classic 1a,2b,3d,4e      1a
2b.3d.e4
   g
(Будь ласка заповнюйте відповідь у вигляді: 'А-1,Б-2,В-3,Г-4')	      )ExamTrainBot.Tests.Questions.FreeQuestion   <text>k__BackingField<points>k__BackingField<answer>k__BackingField<variants>k__BackingFieldrule       Are you a dog?      No
   _
(Будь ласка, будьте уважні при написанні відповіді!)         1   2    3!   5"   7#   78       ,.	
